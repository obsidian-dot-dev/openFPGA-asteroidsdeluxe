module background_lut (
    input wire clk,
    input wire [7:0] index,
    output wire [23:0] pal_rgb_w
);
reg [23:0] pal_rgb;
assign pal_rgb_w = pal_rgb;

always @(posedge clk) begin
  case(index)
    8'd0 : pal_rgb <= 24'h000000;
    8'd1 : pal_rgb <= 24'h030005;
    8'd2 : pal_rgb <= 24'h000306;
    8'd3 : pal_rgb <= 24'h02030f;
    8'd4 : pal_rgb <= 24'h090301;
    8'd5 : pal_rgb <= 24'h050516;
    8'd6 : pal_rgb <= 24'h110513;
    8'd7 : pal_rgb <= 24'h13070f;
    8'd8 : pal_rgb <= 24'h080a1e;
    8'd9 : pal_rgb <= 24'h16090a;
    8'd10 : pal_rgb <= 24'h010f1c;
    8'd11 : pal_rgb <= 24'h03110a;
    8'd12 : pal_rgb <= 24'h120e04;
    8'd13 : pal_rgb <= 24'h1c0b0e;
    8'd14 : pal_rgb <= 24'h240a12;
    8'd15 : pal_rgb <= 24'h1b0d14;
    8'd16 : pal_rgb <= 24'h04161a;
    8'd17 : pal_rgb <= 24'h061803;
    8'd18 : pal_rgb <= 24'h0b142d;
    8'd19 : pal_rgb <= 24'h121231;
    8'd20 : pal_rgb <= 24'h191039;
    8'd21 : pal_rgb <= 24'h1a1506;
    8'd22 : pal_rgb <= 24'h021c14;
    8'd23 : pal_rgb <= 24'h251025;
    8'd24 : pal_rgb <= 24'h19151e;
    8'd25 : pal_rgb <= 24'h151627;
    8'd26 : pal_rgb <= 24'h1f1327;
    8'd27 : pal_rgb <= 24'h0a1a27;
    8'd28 : pal_rgb <= 24'h0c1d01;
    8'd29 : pal_rgb <= 24'h1e1803;
    8'd30 : pal_rgb <= 24'h192139;
    8'd31 : pal_rgb <= 24'h1e2132;
    8'd32 : pal_rgb <= 24'h241f37;
    8'd33 : pal_rgb <= 24'h22212c;
    8'd34 : pal_rgb <= 24'h0a2d13;
    8'd35 : pal_rgb <= 24'h033105;
    8'd36 : pal_rgb <= 24'h0a2d22;
    8'd37 : pal_rgb <= 24'h282513;
    8'd38 : pal_rgb <= 24'h122938;
    8'd39 : pal_rgb <= 24'h072d33;
    8'd40 : pal_rgb <= 24'h182931;
    8'd41 : pal_rgb <= 24'h2f2325;
    8'd42 : pal_rgb <= 24'h242448;
    8'd43 : pal_rgb <= 24'h2e223d;
    8'd44 : pal_rgb <= 24'h27271c;
    8'd45 : pal_rgb <= 24'h2b224e;
    8'd46 : pal_rgb <= 24'h3a2124;
    8'd47 : pal_rgb <= 24'h282908;
    8'd48 : pal_rgb <= 24'h1d2d06;
    8'd49 : pal_rgb <= 24'h352232;
    8'd50 : pal_rgb <= 24'h1d2848;
    8'd51 : pal_rgb <= 24'h262827;
    8'd52 : pal_rgb <= 24'h242c44;
    8'd53 : pal_rgb <= 24'h2f2943;
    8'd54 : pal_rgb <= 24'h282c3d;
    8'd55 : pal_rgb <= 24'h2d2c36;
    8'd56 : pal_rgb <= 24'h313655;
    8'd57 : pal_rgb <= 24'h2f365d;
    8'd58 : pal_rgb <= 24'h124703;
    8'd59 : pal_rgb <= 24'h303849;
    8'd60 : pal_rgb <= 24'h3a3549;
    8'd61 : pal_rgb <= 24'h383838;
    8'd62 : pal_rgb <= 24'h0d4729;
    8'd63 : pal_rgb <= 24'h0e463a;
    8'd64 : pal_rgb <= 24'h0e4917;
    8'd65 : pal_rgb <= 24'h7d261f;
    8'd66 : pal_rgb <= 24'h164347;
    8'd67 : pal_rgb <= 24'h403c16;
    8'd68 : pal_rgb <= 24'h433843;
    8'd69 : pal_rgb <= 24'h3f376c;
    8'd70 : pal_rgb <= 24'h334217;
    8'd71 : pal_rgb <= 24'h40385e;
    8'd72 : pal_rgb <= 24'h23443c;
    8'd73 : pal_rgb <= 24'h2b404e;
    8'd74 : pal_rgb <= 24'h2b405b;
    8'd75 : pal_rgb <= 24'h28452b;
    8'd76 : pal_rgb <= 24'h35412b;
    8'd77 : pal_rgb <= 24'h3b3d45;
    8'd78 : pal_rgb <= 24'h2f4145;
    8'd79 : pal_rgb <= 24'h035407;
    8'd80 : pal_rgb <= 24'h403e2d;
    8'd81 : pal_rgb <= 24'h384406;
    8'd82 : pal_rgb <= 24'h493a3e;
    8'd83 : pal_rgb <= 24'h33413d;
    8'd84 : pal_rgb <= 24'h4e3a2e;
    8'd85 : pal_rgb <= 24'h3a4169;
    8'd86 : pal_rgb <= 24'h3e4262;
    8'd87 : pal_rgb <= 24'h3c4456;
    8'd88 : pal_rgb <= 24'h464156;
    8'd89 : pal_rgb <= 24'h444443;
    8'd90 : pal_rgb <= 24'h14622a;
    8'd91 : pal_rgb <= 24'h106615;
    8'd92 : pal_rgb <= 24'h5f4762;
    8'd93 : pal_rgb <= 24'h4a4d6e;
    8'd94 : pal_rgb <= 24'h16623e;
    8'd95 : pal_rgb <= 24'h415261;
    8'd96 : pal_rgb <= 24'h4e4e65;
    8'd97 : pal_rgb <= 24'h514e5d;
    8'd98 : pal_rgb <= 24'h564e4f;
    8'd99 : pal_rgb <= 24'h215f50;
    8'd100 : pal_rgb <= 24'h544c83;
    8'd101 : pal_rgb <= 24'h326015;
    8'd102 : pal_rgb <= 24'h126c00;
    8'd103 : pal_rgb <= 24'h315f2d;
    8'd104 : pal_rgb <= 24'h744c1b;
    8'd105 : pal_rgb <= 24'h2f5f41;
    8'd106 : pal_rgb <= 24'h315c5e;
    8'd107 : pal_rgb <= 24'h405671;
    8'd108 : pal_rgb <= 24'h6a4c53;
    8'd109 : pal_rgb <= 24'h4d5b17;
    8'd110 : pal_rgb <= 24'h5a4f76;
    8'd111 : pal_rgb <= 24'h654f53;
    8'd112 : pal_rgb <= 24'h385d53;
    8'd113 : pal_rgb <= 24'h425d41;
    8'd114 : pal_rgb <= 24'h685145;
    8'd115 : pal_rgb <= 24'h4b585e;
    8'd116 : pal_rgb <= 24'h58545e;
    8'd117 : pal_rgb <= 24'h4b5c30;
    8'd118 : pal_rgb <= 24'h5c5731;
    8'd119 : pal_rgb <= 24'h595744;
    8'd120 : pal_rgb <= 24'h555755;
    8'd121 : pal_rgb <= 24'h4c5a55;
    8'd122 : pal_rgb <= 24'h4e5b43;
    8'd123 : pal_rgb <= 24'h6b526e;
    8'd124 : pal_rgb <= 24'h4c5d6d;
    8'd125 : pal_rgb <= 24'h565979;
    8'd126 : pal_rgb <= 24'h5b5968;
    8'd127 : pal_rgb <= 24'h595971;
    8'd128 : pal_rgb <= 24'h61595b;
    8'd129 : pal_rgb <= 24'h178017;
    8'd130 : pal_rgb <= 24'h1b7d2e;
    8'd131 : pal_rgb <= 24'h5a6780;
    8'd132 : pal_rgb <= 24'h4a6d77;
    8'd133 : pal_rgb <= 24'h357c1a;
    8'd134 : pal_rgb <= 24'h63686d;
    8'd135 : pal_rgb <= 24'h666865;
    8'd136 : pal_rgb <= 24'h2c7c59;
    8'd137 : pal_rgb <= 24'h2f7d45;
    8'd138 : pal_rgb <= 24'h6a6681;
    8'd139 : pal_rgb <= 24'h3a7c32;
    8'd140 : pal_rgb <= 24'h7c6186;
    8'd141 : pal_rgb <= 24'h3b7868;
    8'd142 : pal_rgb <= 24'h935e5a;
    8'd143 : pal_rgb <= 24'h6e6593;
    8'd144 : pal_rgb <= 24'h5e6d7b;
    8'd145 : pal_rgb <= 24'h796485;
    8'd146 : pal_rgb <= 24'h4f746a;
    8'd147 : pal_rgb <= 24'h5b706e;
    8'd148 : pal_rgb <= 24'h4a794a;
    8'd149 : pal_rgb <= 24'h7a6865;
    8'd150 : pal_rgb <= 24'h437a5b;
    8'd151 : pal_rgb <= 24'h59754a;
    8'd152 : pal_rgb <= 24'h7e685c;
    8'd153 : pal_rgb <= 24'h796b4b;
    8'd154 : pal_rgb <= 24'h77696f;
    8'd155 : pal_rgb <= 24'h6a6c7d;
    8'd156 : pal_rgb <= 24'h617165;
    8'd157 : pal_rgb <= 24'h57755b;
    8'd158 : pal_rgb <= 24'h6a723c;
    8'd159 : pal_rgb <= 24'h58792e;
    8'd160 : pal_rgb <= 24'h67724b;
    8'd161 : pal_rgb <= 24'h6c732f;
    8'd162 : pal_rgb <= 24'h64725b;
    8'd163 : pal_rgb <= 24'h736b7c;
    8'd164 : pal_rgb <= 24'h567a3e;
    8'd165 : pal_rgb <= 24'h6f6f67;
    8'd166 : pal_rgb <= 24'h72705f;
    8'd167 : pal_rgb <= 24'hab6156;
    8'd168 : pal_rgb <= 24'h84723b;
    8'd169 : pal_rgb <= 24'h737572;
    8'd170 : pal_rgb <= 24'h71757a;
    8'd171 : pal_rgb <= 24'ha16c53;
    8'd172 : pal_rgb <= 24'ha37046;
    8'd173 : pal_rgb <= 24'h31982a;
    8'd174 : pal_rgb <= 24'h2b9c16;
    8'd175 : pal_rgb <= 24'h9a7656;
    8'd176 : pal_rgb <= 24'h279b47;
    8'd177 : pal_rgb <= 24'h6b8929;
    8'd178 : pal_rgb <= 24'h319759;
    8'd179 : pal_rgb <= 24'h439647;
    8'd180 : pal_rgb <= 24'ha1794a;
    8'd181 : pal_rgb <= 24'h41946f;
    8'd182 : pal_rgb <= 24'h4b935a;
    8'd183 : pal_rgb <= 24'h579347;
    8'd184 : pal_rgb <= 24'h808283;
    8'd185 : pal_rgb <= 24'h599070;
    8'd186 : pal_rgb <= 24'h71887e;
    8'd187 : pal_rgb <= 24'h8d7f82;
    8'd188 : pal_rgb <= 24'h858932;
    8'd189 : pal_rgb <= 24'h579736;
    8'd190 : pal_rgb <= 24'h84847c;
    8'd191 : pal_rgb <= 24'h669252;
    8'd192 : pal_rgb <= 24'h6e8d72;
    8'd193 : pal_rgb <= 24'h928462;
    8'd194 : pal_rgb <= 24'h629361;
    8'd195 : pal_rgb <= 24'h888675;
    8'd196 : pal_rgb <= 24'h968273;
    8'd197 : pal_rgb <= 24'h758f53;
    8'd198 : pal_rgb <= 24'h7d8a73;
    8'd199 : pal_rgb <= 24'h728f62;
    8'd200 : pal_rgb <= 24'h6b9546;
    8'd201 : pal_rgb <= 24'h8b886f;
    8'd202 : pal_rgb <= 24'h858d55;
    8'd203 : pal_rgb <= 24'h878e47;
    8'd204 : pal_rgb <= 24'h7b9247;
    8'd205 : pal_rgb <= 24'h828e65;
    8'd206 : pal_rgb <= 24'h8c8b66;
    8'd207 : pal_rgb <= 24'ha08a42;
    8'd208 : pal_rgb <= 24'ha18e54;
    8'd209 : pal_rgb <= 24'h45af3b;
    8'd210 : pal_rgb <= 24'h42b327;
    8'd211 : pal_rgb <= 24'h4aac65;
    8'd212 : pal_rgb <= 24'h44b054;
    8'd213 : pal_rgb <= 24'h9f9370;
    8'd214 : pal_rgb <= 24'h61a86f;
    8'd215 : pal_rgb <= 24'ha49566;
    8'd216 : pal_rgb <= 24'h63ad40;
    8'd217 : pal_rgb <= 24'h989d45;
    8'd218 : pal_rgb <= 24'h73aa43;
    8'd219 : pal_rgb <= 24'h5eaf57;
    8'd220 : pal_rgb <= 24'h6faa55;
    8'd221 : pal_rgb <= 24'h68ac66;
    8'd222 : pal_rgb <= 24'h91a345;
    8'd223 : pal_rgb <= 24'h82a844;
    8'd224 : pal_rgb <= 24'haa9687;
    8'd225 : pal_rgb <= 24'h979e87;
    8'd226 : pal_rgb <= 24'ha09f5b;
    8'd227 : pal_rgb <= 24'h81aa59;
    8'd228 : pal_rgb <= 24'h7aaa76;
    8'd229 : pal_rgb <= 24'ha09f79;
    8'd230 : pal_rgb <= 24'h7fab6a;
    8'd231 : pal_rgb <= 24'h9fa26a;
    8'd232 : pal_rgb <= 24'h91a85c;
    8'd233 : pal_rgb <= 24'h98a47a;
    8'd234 : pal_rgb <= 24'ha39f8d;
    8'd235 : pal_rgb <= 24'h8cab8a;
    8'd236 : pal_rgb <= 24'h92ac6f;
    8'd237 : pal_rgb <= 24'h8fac7d;
    8'd238 : pal_rgb <= 24'ha5a8a3;
    8'd239 : pal_rgb <= 24'ha1ab94;
    8'd240 : pal_rgb <= 24'h5fc73d;
    8'd241 : pal_rgb <= 24'h5ec566;
    8'd242 : pal_rgb <= 24'h61c653;
    8'd243 : pal_rgb <= 24'h7ec54a;
    8'd244 : pal_rgb <= 24'h81c541;
    8'd245 : pal_rgb <= 24'h79c65a;
    8'd246 : pal_rgb <= 24'h76c66b;
    8'd247 : pal_rgb <= 24'h7dc47c;
    8'd248 : pal_rgb <= 24'h8dc558;
    8'd249 : pal_rgb <= 24'h87c571;
    8'd250 : pal_rgb <= 24'h9dc45e;
    8'd251 : pal_rgb <= 24'h95c687;
    8'd252 : pal_rgb <= 24'ha2c675;
    8'd253 : pal_rgb <= 24'hbac0b9;
    8'd254 : pal_rgb <= 24'hb7c499;
    8'd255 : pal_rgb <= 24'hb8c4ad;
  endcase
end

endmodule