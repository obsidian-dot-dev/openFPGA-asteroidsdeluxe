//
// User core top-level
//
// Instantiated by the real top-level: apf_top
//

`default_nettype none

module core_top (

//
// physical connections
//

///////////////////////////////////////////////////
// clock inputs 74.25mhz. not phase aligned, so treat these domains as asynchronous

input   wire            clk_74a, // mainclk1
input   wire            clk_74b, // mainclk1 

///////////////////////////////////////////////////
// cartridge interface
// switches between 3.3v and 5v mechanically
// output enable for multibit translators controlled by pic32

// GBA AD[15:8]
inout   wire    [7:0]   cart_tran_bank2,
output  wire            cart_tran_bank2_dir,

// GBA AD[7:0]
inout   wire    [7:0]   cart_tran_bank3,
output  wire            cart_tran_bank3_dir,

// GBA A[23:16]
inout   wire    [7:0]   cart_tran_bank1,
output  wire            cart_tran_bank1_dir,

// GBA [7] PHI#
// GBA [6] WR#
// GBA [5] RD#
// GBA [4] CS1#/CS#
//     [3:0] unwired
inout   wire    [7:4]   cart_tran_bank0,
output  wire            cart_tran_bank0_dir,

// GBA CS2#/RES#
inout   wire            cart_tran_pin30,
output  wire            cart_tran_pin30_dir,
// when GBC cart is inserted, this signal when low or weak will pull GBC /RES low with a special circuit
// the goal is that when unconfigured, the FPGA weak pullups won't interfere.
// thus, if GBC cart is inserted, FPGA must drive this high in order to let the level translators
// and general IO drive this pin.
output  wire            cart_pin30_pwroff_reset,

// GBA IRQ/DRQ
inout   wire            cart_tran_pin31,
output  wire            cart_tran_pin31_dir,

// infrared
input   wire            port_ir_rx,
output  wire            port_ir_tx,
output  wire            port_ir_rx_disable, 

// GBA link port
inout   wire            port_tran_si,
output  wire            port_tran_si_dir,
inout   wire            port_tran_so,
output  wire            port_tran_so_dir,
inout   wire            port_tran_sck,
output  wire            port_tran_sck_dir,
inout   wire            port_tran_sd,
output  wire            port_tran_sd_dir,
 
///////////////////////////////////////////////////
// cellular psram 0 and 1, two chips (64mbit x2 dual die per chip)

output  wire    [21:16] cram0_a,
inout   wire    [15:0]  cram0_dq,
input   wire            cram0_wait,
output  wire            cram0_clk,
output  wire            cram0_adv_n,
output  wire            cram0_cre,
output  wire            cram0_ce0_n,
output  wire            cram0_ce1_n,
output  wire            cram0_oe_n,
output  wire            cram0_we_n,
output  wire            cram0_ub_n,
output  wire            cram0_lb_n,

output  wire    [21:16] cram1_a,
inout   wire    [15:0]  cram1_dq,
input   wire            cram1_wait,
output  wire            cram1_clk,
output  wire            cram1_adv_n,
output  wire            cram1_cre,
output  wire            cram1_ce0_n,
output  wire            cram1_ce1_n,
output  wire            cram1_oe_n,
output  wire            cram1_we_n,
output  wire            cram1_ub_n,
output  wire            cram1_lb_n,

///////////////////////////////////////////////////
// sdram, 512mbit 16bit

output  wire    [12:0]  dram_a,
output  wire    [1:0]   dram_ba,
inout   wire    [15:0]  dram_dq,
output  wire    [1:0]   dram_dqm,
output  wire            dram_clk,
output  wire            dram_cke,
output  wire            dram_ras_n,
output  wire            dram_cas_n,
output  wire            dram_we_n,

///////////////////////////////////////////////////
// sram, 1mbit 16bit

output  wire    [16:0]  sram_a,
inout   wire    [15:0]  sram_dq,
output  wire            sram_oe_n,
output  wire            sram_we_n,
output  wire            sram_ub_n,
output  wire            sram_lb_n,

///////////////////////////////////////////////////
// vblank driven by dock for sync in a certain mode

input   wire            vblank,

///////////////////////////////////////////////////
// i/o to 6515D breakout usb uart

output  wire            dbg_tx,
input   wire            dbg_rx,

///////////////////////////////////////////////////
// i/o pads near jtag connector user can solder to

output  wire            user1,
input   wire            user2,

///////////////////////////////////////////////////
// RFU internal i2c bus 

inout   wire            aux_sda,
output  wire            aux_scl,

///////////////////////////////////////////////////
// RFU, do not use
output  wire            vpll_feed,


//
// logical connections
//

///////////////////////////////////////////////////
// video, audio output to scaler
output  wire    [23:0]  video_rgb,
output  wire            video_rgb_clock,
output  wire            video_rgb_clock_90,
output  wire            video_de,
output  wire            video_skip,
output  wire            video_vs,
output  wire            video_hs,
    
output  wire            audio_mclk,
input   wire            audio_adc,
output  wire            audio_dac,
output  wire            audio_lrck,

///////////////////////////////////////////////////
// bridge bus connection
// synchronous to clk_74a
output  wire            bridge_endian_little,
input   wire    [31:0]  bridge_addr,
input   wire            bridge_rd,
output  reg     [31:0]  bridge_rd_data,
input   wire            bridge_wr,
input   wire    [31:0]  bridge_wr_data,

///////////////////////////////////////////////////
// controller data
// 
// key bitmap:
//   [0]    dpad_up
//   [1]    dpad_down
//   [2]    dpad_left
//   [3]    dpad_right
//   [4]    face_a
//   [5]    face_b
//   [6]    face_x
//   [7]    face_y
//   [8]    trig_l1
//   [9]    trig_r1
//   [10]   trig_l2
//   [11]   trig_r2
//   [12]   trig_l3
//   [13]   trig_r3
//   [14]   face_select
//   [15]   face_start
// joy values - unsigned
//   [ 7: 0] lstick_x
//   [15: 8] lstick_y
//   [23:16] rstick_x
//   [31:24] rstick_y
// trigger values - unsigned
//   [ 7: 0] ltrig
//   [15: 8] rtrig
//
input   wire    [31:0]  cont1_key,
input   wire    [31:0]  cont2_key,
input   wire    [31:0]  cont3_key,
input   wire    [31:0]  cont4_key,
input   wire    [31:0]  cont1_joy,
input   wire    [31:0]  cont2_joy,
input   wire    [31:0]  cont3_joy,
input   wire    [31:0]  cont4_joy,
input   wire    [15:0]  cont1_trig,
input   wire    [15:0]  cont2_trig,
input   wire    [15:0]  cont3_trig,
input   wire    [15:0]  cont4_trig
    
);

// not using the IR port, so turn off both the LED, and
// disable the receive circuit to save power
assign port_ir_tx = 0;
assign port_ir_rx_disable = 1;

// bridge endianness
assign bridge_endian_little = 0;

// cart is unused, so set all level translators accordingly
// directions are 0:IN, 1:OUT
assign cart_tran_bank3 = 8'hzz;
assign cart_tran_bank3_dir = 1'b0;
assign cart_tran_bank2 = 8'hzz;
assign cart_tran_bank2_dir = 1'b0;
assign cart_tran_bank1 = 8'hzz;
assign cart_tran_bank1_dir = 1'b0;
assign cart_tran_bank0 = 4'hf;
assign cart_tran_bank0_dir = 1'b1;
assign cart_tran_pin30 = 1'b0;      // reset or cs2, we let the hw control it by itself
assign cart_tran_pin30_dir = 1'bz;
assign cart_pin30_pwroff_reset = 1'b0;  // hardware can control this
assign cart_tran_pin31 = 1'bz;      // input
assign cart_tran_pin31_dir = 1'b0;  // input

// link port is input only
assign port_tran_so = 1'bz;
assign port_tran_so_dir = 1'b0;     // SO is output only
assign port_tran_si = 1'bz;
assign port_tran_si_dir = 1'b0;     // SI is input only
assign port_tran_sck = 1'bz;
assign port_tran_sck_dir = 1'b0;    // clock direction can change
assign port_tran_sd = 1'bz;
assign port_tran_sd_dir = 1'b0;     // SD is input and not used

// tie off the rest of the pins we are not using
assign cram0_a = 'h0;
assign cram0_dq = {16{1'bZ}};
assign cram0_clk = 0;
assign cram0_adv_n = 1;
assign cram0_cre = 0;
assign cram0_ce0_n = 1;
assign cram0_ce1_n = 1;
assign cram0_oe_n = 1;
assign cram0_we_n = 1;
assign cram0_ub_n = 1;
assign cram0_lb_n = 1;

assign cram1_a = 'h0;
assign cram1_dq = {16{1'bZ}};
assign cram1_clk = 0;
assign cram1_adv_n = 1;
assign cram1_cre = 0;
assign cram1_ce0_n = 1;
assign cram1_ce1_n = 1;
assign cram1_oe_n = 1;
assign cram1_we_n = 1;
assign cram1_ub_n = 1;
assign cram1_lb_n = 1;

assign dram_a = 'h0;
assign dram_ba = 'h0;
assign dram_dq = {16{1'bZ}};
assign dram_dqm = 'h0;
assign dram_clk = 'h0;
assign dram_cke = 'h0;
assign dram_ras_n = 'h1;
assign dram_cas_n = 'h1;
assign dram_we_n = 'h1;

// assign sram_a = 'h0;
// assign sram_dq = {16{1'bZ}};
// assign sram_oe_n  = 1;
// assign sram_we_n  = 1;
// assign sram_ub_n  = 1;
// assign sram_lb_n  = 1;

assign dbg_tx = 1'bZ;
assign user1 = 1'bZ;
assign aux_scl = 1'bZ;
assign vpll_feed = 1'bZ;


// for bridge write data, we just broadcast it to all bus devices
// for bridge read data, we have to mux it
// add your own devices here
always @(*) begin
    casex(bridge_addr)
    default: begin
        bridge_rd_data <= 0;
    end
    32'h10xxxxxx: begin
        // example
        // bridge_rd_data <= example_device_data;
        bridge_rd_data <= 0;
    end
    32'hF8xxxxxx: begin
        bridge_rd_data <= cmd_bridge_rd_data;
    end
    endcase
end


//
// host/target command handler
//
    wire            reset_n;                // driven by host commands, can be used as core-wide reset
    wire    [31:0]  cmd_bridge_rd_data;
    
// bridge host commands
// synchronous to clk_74a
    wire            status_boot_done = pll_core_locked; 
    wire            status_setup_done = pll_core_locked; // rising edge triggers a target command
    wire            status_running = reset_n; // we are running as soon as reset_n goes high

    wire            dataslot_requestread;
    wire    [15:0]  dataslot_requestread_id;
    wire            dataslot_requestread_ack = 1;
    wire            dataslot_requestread_ok = 1;

    wire            dataslot_requestwrite;
    wire    [15:0]  dataslot_requestwrite_id;
    wire            dataslot_requestwrite_ack = 1;
    wire            dataslot_requestwrite_ok = 1;

    wire            dataslot_allcomplete;

    wire            savestate_supported;
    wire    [31:0]  savestate_addr;
    wire    [31:0]  savestate_size;
    wire    [31:0]  savestate_maxloadsize;

    wire            savestate_start;
    wire            savestate_start_ack;
    wire            savestate_start_busy;
    wire            savestate_start_ok;
    wire            savestate_start_err;

    wire            savestate_load;
    wire            savestate_load_ack;
    wire            savestate_load_busy;
    wire            savestate_load_ok;
    wire            savestate_load_err;
    
    wire            osnotify_inmenu;

// bridge target commands
// synchronous to clk_74a


// bridge data slot access

    wire    [9:0]   datatable_addr;
    wire            datatable_wren;
    wire    [31:0]  datatable_data;
    wire    [31:0]  datatable_q;

core_bridge_cmd icb (

    .clk                ( clk_74a ),
    .reset_n            ( reset_n ),

    .bridge_endian_little   ( bridge_endian_little ),
    .bridge_addr            ( bridge_addr ),
    .bridge_rd              ( bridge_rd ),
    .bridge_rd_data         ( cmd_bridge_rd_data ),
    .bridge_wr              ( bridge_wr ),
    .bridge_wr_data         ( bridge_wr_data ),
    
    .status_boot_done       ( status_boot_done ),
    .status_setup_done      ( status_setup_done ),
    .status_running         ( status_running ),

    .dataslot_requestread       ( dataslot_requestread ),
    .dataslot_requestread_id    ( dataslot_requestread_id ),
    .dataslot_requestread_ack   ( dataslot_requestread_ack ),
    .dataslot_requestread_ok    ( dataslot_requestread_ok ),

    .dataslot_requestwrite      ( dataslot_requestwrite ),
    .dataslot_requestwrite_id   ( dataslot_requestwrite_id ),
    .dataslot_requestwrite_ack  ( dataslot_requestwrite_ack ),
    .dataslot_requestwrite_ok   ( dataslot_requestwrite_ok ),

    .dataslot_allcomplete   ( dataslot_allcomplete ),

    .savestate_supported    ( savestate_supported ),
    .savestate_addr         ( savestate_addr ),
    .savestate_size         ( savestate_size ),
    .savestate_maxloadsize  ( savestate_maxloadsize ),

    .savestate_start        ( savestate_start ),
    .savestate_start_ack    ( savestate_start_ack ),
    .savestate_start_busy   ( savestate_start_busy ),
    .savestate_start_ok     ( savestate_start_ok ),
    .savestate_start_err    ( savestate_start_err ),

    .savestate_load         ( savestate_load ),
    .savestate_load_ack     ( savestate_load_ack ),
    .savestate_load_busy    ( savestate_load_busy ),
    .savestate_load_ok      ( savestate_load_ok ),
    .savestate_load_err     ( savestate_load_err ),

    .osnotify_inmenu        ( osnotify_inmenu ),
    
    .datatable_addr         ( datatable_addr ),
    .datatable_wren         ( datatable_wren ),
    .datatable_data         ( datatable_data ),
    .datatable_q            ( datatable_q ),

);



////////////////////////////////////////////////////////////////////////////////////////

wire clk_6;
wire clk_25;
wire clk_25_175;
wire clk_25_175_90deg;
wire clk_50;

wire    pll_core_locked;
    
mf_pllbase mp1 (
    .refclk         ( clk_74a ),
    .rst            ( 0 ),
    
    .outclk_0       ( clk_6 ),
    .outclk_1       ( clk_25_175_90deg ),
    .outclk_2       ( clk_50 ),
    .outclk_3       ( clk_25 ),
    .outclk_4       ( clk_25_175 ),

    .locked         ( pll_core_locked )
);

///////////////////////////////////////////////
// Core Settings
///////////////////////////////////////////////

reg [1:0] cs_language   = 0;
reg [1:0] cs_ship_count = 0;
reg [1:0] cs_bonus 		= 0;
reg cs_background = 0;
always @(posedge clk_74a) begin
  if(bridge_wr) begin
    casex(bridge_addr)
      32'h80000000: cs_language   <= bridge_wr_data[1:0];
      32'h90000000: cs_ship_count <= bridge_wr_data[1:0];
      32'h10000000: cs_bonus		 <= bridge_wr_data[1:0];
      32'h20000000: cs_background <= bridge_wr_data[0];
    endcase
  end
end

///////////////////////////////////////////////
// Core Audio
///////////////////////////////////////////////

wire [7:0] audio;

sound_i2s #(
    .CHANNEL_WIDTH(8),
    .SIGNED_INPUT (0)
) sound_i2s (
    .clk_74a(clk_74a),
    .clk_audio(clk_6),
    
    .audio_l(audio),
    .audio_r(audio),

    .audio_mclk(audio_mclk),
    .audio_lrck(audio_lrck),
    .audio_dac(audio_dac)
);

///////////////////////////////////////////////
// Core Video
///////////////////////////////////////////////

assign video_rgb_clock = clk_25_175;
assign video_rgb_clock_90 = clk_25_175_90deg;

reg video_de_reg;
reg video_hs_reg;
reg video_vs_reg;
reg [23:0] video_rgb_reg;
reg video_skip_reg;

assign video_de = video_de_reg;
assign video_hs = video_hs_reg;
assign video_vs = video_vs_reg;
assign video_rgb = video_rgb_reg;
assign video_skip = video_skip_reg;

reg hs_prev;
reg vs_prev;
reg de_prev;

always @(posedge clk_25_175) begin
  video_de_reg <= 0;
  video_rgb_reg <= 24'h0;

  if (~(vblank_asteroids || hblank)) begin
    video_de_reg <= 1;

	 if (cs_background && !r2 && !g2 && !b2) begin
     video_rgb_reg[23:16] <= {2'b0, pal_rgb_w[23:18]};
     video_rgb_reg[15:8] <= {2'b0, pal_rgb_w[15:10]};
     video_rgb_reg[7:0] <= {2'b0, pal_rgb_w[7:2]};
	 end
	 else begin
		 video_rgb_reg[23:16] <= {2{r2}};
		 video_rgb_reg[15:8]  <= {2{g2}};
		 video_rgb_reg[7:0]   <= {2{b2}};
	 end
  end

  video_hs_reg <= ~hs_prev && hs;
  video_vs_reg <= ~vs_prev && vs;
  hs_prev <= hs;
  vs_prev <= vs;
end

///////////////////////////////////////////////
// Background
///////////////////////////////////////////////

reg [18:0] bg_addr;
reg [18:0] bg_base_addr;

reg [8:0] bg_row;
wire [7:0] bg_pix;

always @(posedge clk_25_175) begin
  reg vblank_prev;
  reg hblank_prev; 
  vblank_prev <= vblank_asteroids;
  hblank_prev <= hblank;
  if (vblank_asteroids) begin
    bg_base_addr <= 0;
    bg_addr <= 2;
	  bg_row <= 0;
  end  
  if (!vblank_asteroids && !hblank) begin
    if (!vblank_asteroids && vblank_prev) begin
	   bg_base_addr <= 2;
		 bg_row <= 0;
	 end
	 else if (hblank_prev && !hblank) begin
	   if (bg_row != 0) begin
        bg_base_addr <= bg_base_addr + 19'd640;
		  bg_addr <= bg_base_addr + 19'd640;
		  bg_row <= bg_row + 9'd1;
		end
		else begin
		  bg_base_addr <= bg_base_addr + 19'd640;
		  bg_addr <= bg_base_addr + 19'd640;
		end
	 end
	 else if (!hblank_prev && !hblank) begin
		bg_addr <= bg_addr + 19'd1;
	 end
  end
end

reg [7:0] bg_bram_pix;

// Lower 64KB stored in bram
wire bg_bram_download;
assign bg_bram_download = (ioctl_wr && ioctl_addr[24] == 1 && ioctl_addr[18:16] == 0);

// Upper 256KB stored in sram
wire bg_sram_download;
assign bg_sram_download = (ioctl_wr && ioctl_addr[24] == 1 && ioctl_addr[18:16] != 3'b0);

wire [15:0] bg_sram_load;
reg [15:0] bg_sram_store;
reg [7:0]  bg_low;
reg [16:0] bg_sram_addr;
reg [7:0]  bg_sram_pix;

wire [2:0] ioctl_bank;
wire [2:0] bg_sram_bank;

assign ioctl_bank = ioctl_addr[18:16] - 3'b1;
assign bg_sram_bank = bg_addr[18:16] - 3'b1;

reg bg_sram_wren;

// Remaining chunk of background data is in SRAM.
always @(posedge clk_50) begin
  // If downloading the image data...
  if (bg_sram_download) begin
     if (ioctl_addr[0] == 0) begin
	   bg_low <= ioctl_dout;
	 end
	 else if (ioctl_addr[0] == 1) begin
	   bg_sram_store[15:8] <= ioctl_dout;
		 bg_sram_store[7:0] <= bg_low;
		 bg_sram_addr <= {ioctl_bank[1:0], ioctl_addr[15:1]}; // account for the 64K offset
	 end
  end
  // If reading the image data back...
  else begin
    bg_sram_addr <= {bg_sram_bank[1:0], bg_addr[15:1]}; // account for the 64K offset
    if (bg_addr[0] == 0) begin
	   bg_sram_pix <= bg_sram_load[15:8];
	 end
    else begin
	   bg_sram_pix <= bg_sram_load[7:0];
	 end
  end
end

assign bg_pix = bg_addr[18:16] == 0 ? bg_bram_pix : bg_sram_pix;

// 1st chunk of background data is in DPRAM.
dpram #(
  .addr_width_g(16),  // 64 KB
  .data_width_g(8),
  .num_words_g(65536)
) bg_bram1 (
  .address_a(ioctl_addr[15:0]),
  .address_b(bg_addr[15:0]),
  .clock_a(clk_50),
  .clock_b(clk_50),
  .data_a(ioctl_dout),
  .enable_a(1'b1),
  .enable_b(1'b1),
  .wren_a(bg_bram_download),
  .wren_b(1'b0),
  .q_b(bg_bram_pix),
);

// Remaining background image data is stored in SRAM.
sram_storage sram_storage(
	.wr_en(bg_sram_download),
	
	.addr(bg_sram_addr),
	.din(bg_sram_store),
	.dout(bg_sram_load),
	
	.sram_a(sram_a),
	.sram_dq(sram_dq),
	.sram_oe_n(sram_oe_n),
	.sram_we_n(sram_we_n),
	.sram_ub_n(sram_ub_n),
	.sram_lb_n(sram_lb_n),
);

// Background image is 8bpp, indexed.  We need a lut
// to convert the index values to 24-bit RGB data.
wire [23:0] pal_rgb_w;

background_lut background_lut(
  .clk(clk_50),
  .index(bg_pix),
  .pal_rgb_w(pal_rgb_w),
);


///////////////////////////////////////////////
// Core Instance
///////////////////////////////////////////////

wire        ioctl_wr;
wire [24:0] ioctl_addr;
wire  [7:0] ioctl_dout;

data_loader #(
    .WRITE_MEM_CLOCK_DELAY(4)
) rom_loader (
    .clk_74a(clk_74a),
    .clk_memory(clk_25),

    .bridge_wr(bridge_wr),
    .bridge_endian_little(bridge_endian_little),
    .bridge_addr(bridge_addr),
    .bridge_wr_data(bridge_wr_data),

    .write_en(ioctl_wr),
    .write_addr(ioctl_addr),
    .write_data(ioctl_dout)
);

wire [31:0] cont1_key_s;
wire [31:0] cont2_key_s;

synch_2 #(
  .WIDTH(32)
) cont1_s (
  cont1_key,
  cont1_key_s,
  clk_6
);

synch_2 #(
  .WIDTH(32)
) cont2_s (
  cont2_key,
  cont2_key_s,
  clk_6
);

wire [7:0] BUTTON = {
    ~(cont1_key_s[3] | cont2_key_s[3]),  // right
    ~(cont1_key_s[2] | cont2_key_s[2]),  // left
    ~cont1_key_s[15],                    // P1 Start
    ~cont2_key_s[15],                    // P2 Start
    ~(cont1_key_s[4] | cont2_key_s[4]),  // fire
    ~(cont1_key_s[7] | cont2_key_s[7]),  // ???
    ~(cont1_key_s[6] | cont2_key_s[6]),  // thrust
    ~(cont1_key_s[5] | cont2_key_s[5])   // hyperspace
};

wire hblank, vblank_asteroids;
wire hs, vs;
wire [3:0] r,g,b;

reg [3:0] r2;
reg [3:0] g2;
reg [3:0] b2;

always @(posedge clk_50) begin
  r2 <= r;
  g2 <= g;
  b2 <= b;
end

ASTEROIDS_TOP ASTEROIDS_TOP
(
	.dn_addr(ioctl_addr[15:0]),
	.dn_data(ioctl_dout),
	.dn_wr(ioctl_wr && (ioctl_addr[24] == 0)),	
	.clk_6(clk_6),
	.clk_25(clk_25),

	.BUTTON(BUTTON),
	.BONUS(cs_bonus),
//	--.SELF_TEST_SWITCH_L(~cs_bonus), 
	.LANG(cs_language),
	.SHIPS(cs_ship_count),
	.AUDIO_OUT(audio),
  .VIDEO_R_OUT(r),
	.VIDEO_G_OUT(g),
	.VIDEO_B_OUT(b),
	.HSYNC_OUT(hs),
	.VSYNC_OUT(vs),
	.VID_HBLANK(hblank),
	.VID_VBLANK(vblank_asteroids),

	.RESET_L (reset_n),	
);

endmodule
